VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picorv32
  CLASS BLOCK ;
  FOREIGN picorv32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 455.205 BY 465.925 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END clk
  PIN eoi[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END eoi[0]
  PIN eoi[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END eoi[10]
  PIN eoi[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END eoi[11]
  PIN eoi[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END eoi[12]
  PIN eoi[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END eoi[13]
  PIN eoi[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END eoi[14]
  PIN eoi[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END eoi[15]
  PIN eoi[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END eoi[16]
  PIN eoi[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END eoi[17]
  PIN eoi[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END eoi[18]
  PIN eoi[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END eoi[19]
  PIN eoi[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END eoi[1]
  PIN eoi[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END eoi[20]
  PIN eoi[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END eoi[21]
  PIN eoi[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END eoi[22]
  PIN eoi[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END eoi[23]
  PIN eoi[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END eoi[24]
  PIN eoi[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END eoi[25]
  PIN eoi[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END eoi[26]
  PIN eoi[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END eoi[27]
  PIN eoi[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END eoi[28]
  PIN eoi[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END eoi[29]
  PIN eoi[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END eoi[2]
  PIN eoi[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END eoi[30]
  PIN eoi[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END eoi[31]
  PIN eoi[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END eoi[3]
  PIN eoi[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END eoi[4]
  PIN eoi[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END eoi[5]
  PIN eoi[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END eoi[6]
  PIN eoi[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END eoi[7]
  PIN eoi[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END eoi[8]
  PIN eoi[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END eoi[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END irq[15]
  PIN irq[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END irq[16]
  PIN irq[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END irq[17]
  PIN irq[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END irq[18]
  PIN irq[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END irq[19]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END irq[1]
  PIN irq[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END irq[20]
  PIN irq[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END irq[21]
  PIN irq[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END irq[22]
  PIN irq[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END irq[23]
  PIN irq[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END irq[24]
  PIN irq[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END irq[25]
  PIN irq[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END irq[26]
  PIN irq[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END irq[27]
  PIN irq[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END irq[28]
  PIN irq[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END irq[29]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END irq[2]
  PIN irq[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END irq[30]
  PIN irq[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END irq[31]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END irq[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END mem_addr[9]
  PIN mem_instr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END mem_instr
  PIN mem_la_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END mem_la_addr[0]
  PIN mem_la_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END mem_la_addr[10]
  PIN mem_la_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END mem_la_addr[11]
  PIN mem_la_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END mem_la_addr[12]
  PIN mem_la_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END mem_la_addr[13]
  PIN mem_la_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END mem_la_addr[14]
  PIN mem_la_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END mem_la_addr[15]
  PIN mem_la_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END mem_la_addr[16]
  PIN mem_la_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END mem_la_addr[17]
  PIN mem_la_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END mem_la_addr[18]
  PIN mem_la_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END mem_la_addr[19]
  PIN mem_la_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END mem_la_addr[1]
  PIN mem_la_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END mem_la_addr[20]
  PIN mem_la_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END mem_la_addr[21]
  PIN mem_la_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END mem_la_addr[22]
  PIN mem_la_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END mem_la_addr[23]
  PIN mem_la_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END mem_la_addr[24]
  PIN mem_la_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END mem_la_addr[25]
  PIN mem_la_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END mem_la_addr[26]
  PIN mem_la_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END mem_la_addr[27]
  PIN mem_la_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END mem_la_addr[28]
  PIN mem_la_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END mem_la_addr[29]
  PIN mem_la_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END mem_la_addr[2]
  PIN mem_la_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END mem_la_addr[30]
  PIN mem_la_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END mem_la_addr[31]
  PIN mem_la_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END mem_la_addr[3]
  PIN mem_la_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END mem_la_addr[4]
  PIN mem_la_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END mem_la_addr[5]
  PIN mem_la_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END mem_la_addr[6]
  PIN mem_la_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END mem_la_addr[7]
  PIN mem_la_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END mem_la_addr[8]
  PIN mem_la_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END mem_la_addr[9]
  PIN mem_la_read
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END mem_la_read
  PIN mem_la_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END mem_la_wdata[0]
  PIN mem_la_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END mem_la_wdata[10]
  PIN mem_la_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END mem_la_wdata[11]
  PIN mem_la_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END mem_la_wdata[12]
  PIN mem_la_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END mem_la_wdata[13]
  PIN mem_la_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END mem_la_wdata[14]
  PIN mem_la_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END mem_la_wdata[15]
  PIN mem_la_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END mem_la_wdata[16]
  PIN mem_la_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END mem_la_wdata[17]
  PIN mem_la_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END mem_la_wdata[18]
  PIN mem_la_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END mem_la_wdata[19]
  PIN mem_la_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END mem_la_wdata[1]
  PIN mem_la_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END mem_la_wdata[20]
  PIN mem_la_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END mem_la_wdata[21]
  PIN mem_la_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END mem_la_wdata[22]
  PIN mem_la_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END mem_la_wdata[23]
  PIN mem_la_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END mem_la_wdata[24]
  PIN mem_la_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END mem_la_wdata[25]
  PIN mem_la_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END mem_la_wdata[26]
  PIN mem_la_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END mem_la_wdata[27]
  PIN mem_la_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END mem_la_wdata[28]
  PIN mem_la_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END mem_la_wdata[29]
  PIN mem_la_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END mem_la_wdata[2]
  PIN mem_la_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END mem_la_wdata[30]
  PIN mem_la_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END mem_la_wdata[31]
  PIN mem_la_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END mem_la_wdata[3]
  PIN mem_la_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END mem_la_wdata[4]
  PIN mem_la_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END mem_la_wdata[5]
  PIN mem_la_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END mem_la_wdata[6]
  PIN mem_la_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END mem_la_wdata[7]
  PIN mem_la_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END mem_la_wdata[8]
  PIN mem_la_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END mem_la_wdata[9]
  PIN mem_la_write
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END mem_la_write
  PIN mem_la_wstrb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END mem_la_wstrb[0]
  PIN mem_la_wstrb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END mem_la_wstrb[1]
  PIN mem_la_wstrb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END mem_la_wstrb[2]
  PIN mem_la_wstrb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END mem_la_wstrb[3]
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END mem_rdata[9]
  PIN mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END mem_ready
  PIN mem_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END mem_valid
  PIN mem_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END mem_wdata[9]
  PIN mem_wstrb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END mem_wstrb[0]
  PIN mem_wstrb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END mem_wstrb[1]
  PIN mem_wstrb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END mem_wstrb[2]
  PIN mem_wstrb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END mem_wstrb[3]
  PIN pcpi_insn[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END resetn
  PIN trace_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END trace_data[0]
  PIN trace_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END trace_data[10]
  PIN trace_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END trace_data[11]
  PIN trace_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END trace_data[12]
  PIN trace_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END trace_data[13]
  PIN trace_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END trace_data[14]
  PIN trace_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END trace_data[15]
  PIN trace_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END trace_data[16]
  PIN trace_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END trace_data[17]
  PIN trace_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END trace_data[18]
  PIN trace_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END trace_data[19]
  PIN trace_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END trace_data[1]
  PIN trace_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END trace_data[20]
  PIN trace_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END trace_data[21]
  PIN trace_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END trace_data[22]
  PIN trace_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END trace_data[23]
  PIN trace_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END trace_data[24]
  PIN trace_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END trace_data[25]
  PIN trace_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END trace_data[26]
  PIN trace_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END trace_data[27]
  PIN trace_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END trace_data[28]
  PIN trace_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END trace_data[29]
  PIN trace_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END trace_data[2]
  PIN trace_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END trace_data[30]
  PIN trace_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END trace_data[31]
  PIN trace_data[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END trace_data[32]
  PIN trace_data[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END trace_data[33]
  PIN trace_data[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END trace_data[34]
  PIN trace_data[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END trace_data[35]
  PIN trace_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END trace_data[3]
  PIN trace_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END trace_data[4]
  PIN trace_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END trace_data[5]
  PIN trace_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END trace_data[6]
  PIN trace_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END trace_data[7]
  PIN trace_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END trace_data[8]
  PIN trace_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END trace_data[9]
  PIN trace_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END trace_valid
  PIN trap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END trap
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 454.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 454.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 454.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 454.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 454.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 454.480 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 449.610 454.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 449.420 454.325 ;
      LAYER met1 ;
        RECT 5.520 0.380 450.270 454.480 ;
      LAYER met2 ;
        RECT 7.000 4.280 450.240 454.425 ;
        RECT 7.000 0.350 39.370 4.280 ;
        RECT 40.210 0.350 40.290 4.280 ;
        RECT 41.130 0.350 41.210 4.280 ;
        RECT 42.050 0.350 42.130 4.280 ;
        RECT 42.970 0.350 43.050 4.280 ;
        RECT 43.890 0.350 43.970 4.280 ;
        RECT 44.810 0.350 44.890 4.280 ;
        RECT 45.730 0.350 45.810 4.280 ;
        RECT 46.650 0.350 46.730 4.280 ;
        RECT 47.570 0.350 47.650 4.280 ;
        RECT 48.490 0.350 48.570 4.280 ;
        RECT 49.410 0.350 49.490 4.280 ;
        RECT 50.330 0.350 50.410 4.280 ;
        RECT 51.250 0.350 51.330 4.280 ;
        RECT 52.170 0.350 52.250 4.280 ;
        RECT 53.090 0.350 53.170 4.280 ;
        RECT 54.010 0.350 54.090 4.280 ;
        RECT 54.930 0.350 55.010 4.280 ;
        RECT 55.850 0.350 55.930 4.280 ;
        RECT 56.770 0.350 56.850 4.280 ;
        RECT 57.690 0.350 57.770 4.280 ;
        RECT 58.610 0.350 58.690 4.280 ;
        RECT 59.530 0.350 59.610 4.280 ;
        RECT 60.450 0.350 60.530 4.280 ;
        RECT 61.370 0.350 61.450 4.280 ;
        RECT 62.290 0.350 62.370 4.280 ;
        RECT 63.210 0.350 63.290 4.280 ;
        RECT 64.130 0.350 64.210 4.280 ;
        RECT 65.050 0.350 65.130 4.280 ;
        RECT 65.970 0.350 66.050 4.280 ;
        RECT 66.890 0.350 66.970 4.280 ;
        RECT 67.810 0.350 67.890 4.280 ;
        RECT 68.730 0.350 68.810 4.280 ;
        RECT 69.650 0.350 69.730 4.280 ;
        RECT 70.570 0.350 70.650 4.280 ;
        RECT 71.490 0.350 71.570 4.280 ;
        RECT 72.410 0.350 72.490 4.280 ;
        RECT 73.330 0.350 73.410 4.280 ;
        RECT 74.250 0.350 74.330 4.280 ;
        RECT 75.170 0.350 75.250 4.280 ;
        RECT 76.090 0.350 76.170 4.280 ;
        RECT 77.010 0.350 77.090 4.280 ;
        RECT 77.930 0.350 78.010 4.280 ;
        RECT 78.850 0.350 78.930 4.280 ;
        RECT 79.770 0.350 79.850 4.280 ;
        RECT 80.690 0.350 80.770 4.280 ;
        RECT 81.610 0.350 81.690 4.280 ;
        RECT 82.530 0.350 82.610 4.280 ;
        RECT 83.450 0.350 83.530 4.280 ;
        RECT 84.370 0.350 84.450 4.280 ;
        RECT 85.290 0.350 85.370 4.280 ;
        RECT 86.210 0.350 86.290 4.280 ;
        RECT 87.130 0.350 87.210 4.280 ;
        RECT 88.050 0.350 88.130 4.280 ;
        RECT 88.970 0.350 89.050 4.280 ;
        RECT 89.890 0.350 89.970 4.280 ;
        RECT 90.810 0.350 90.890 4.280 ;
        RECT 91.730 0.350 91.810 4.280 ;
        RECT 92.650 0.350 92.730 4.280 ;
        RECT 93.570 0.350 93.650 4.280 ;
        RECT 94.490 0.350 94.570 4.280 ;
        RECT 95.410 0.350 95.490 4.280 ;
        RECT 96.330 0.350 96.410 4.280 ;
        RECT 97.250 0.350 97.330 4.280 ;
        RECT 98.170 0.350 98.250 4.280 ;
        RECT 99.090 0.350 99.170 4.280 ;
        RECT 100.010 0.350 100.090 4.280 ;
        RECT 100.930 0.350 101.010 4.280 ;
        RECT 101.850 0.350 101.930 4.280 ;
        RECT 102.770 0.350 102.850 4.280 ;
        RECT 103.690 0.350 103.770 4.280 ;
        RECT 104.610 0.350 104.690 4.280 ;
        RECT 105.530 0.350 105.610 4.280 ;
        RECT 106.450 0.350 106.530 4.280 ;
        RECT 107.370 0.350 107.450 4.280 ;
        RECT 108.290 0.350 108.370 4.280 ;
        RECT 109.210 0.350 109.290 4.280 ;
        RECT 110.130 0.350 110.210 4.280 ;
        RECT 111.050 0.350 111.130 4.280 ;
        RECT 111.970 0.350 112.050 4.280 ;
        RECT 112.890 0.350 112.970 4.280 ;
        RECT 113.810 0.350 113.890 4.280 ;
        RECT 114.730 0.350 114.810 4.280 ;
        RECT 115.650 0.350 115.730 4.280 ;
        RECT 116.570 0.350 116.650 4.280 ;
        RECT 117.490 0.350 117.570 4.280 ;
        RECT 118.410 0.350 118.490 4.280 ;
        RECT 119.330 0.350 119.410 4.280 ;
        RECT 120.250 0.350 120.330 4.280 ;
        RECT 121.170 0.350 121.250 4.280 ;
        RECT 122.090 0.350 122.170 4.280 ;
        RECT 123.010 0.350 123.090 4.280 ;
        RECT 123.930 0.350 124.010 4.280 ;
        RECT 124.850 0.350 124.930 4.280 ;
        RECT 125.770 0.350 125.850 4.280 ;
        RECT 126.690 0.350 126.770 4.280 ;
        RECT 127.610 0.350 127.690 4.280 ;
        RECT 128.530 0.350 128.610 4.280 ;
        RECT 129.450 0.350 129.530 4.280 ;
        RECT 130.370 0.350 130.450 4.280 ;
        RECT 131.290 0.350 131.370 4.280 ;
        RECT 132.210 0.350 132.290 4.280 ;
        RECT 133.130 0.350 133.210 4.280 ;
        RECT 134.050 0.350 134.130 4.280 ;
        RECT 134.970 0.350 135.050 4.280 ;
        RECT 135.890 0.350 135.970 4.280 ;
        RECT 136.810 0.350 136.890 4.280 ;
        RECT 137.730 0.350 137.810 4.280 ;
        RECT 138.650 0.350 138.730 4.280 ;
        RECT 139.570 0.350 139.650 4.280 ;
        RECT 140.490 0.350 140.570 4.280 ;
        RECT 141.410 0.350 141.490 4.280 ;
        RECT 142.330 0.350 142.410 4.280 ;
        RECT 143.250 0.350 143.330 4.280 ;
        RECT 144.170 0.350 144.250 4.280 ;
        RECT 145.090 0.350 145.170 4.280 ;
        RECT 146.010 0.350 146.090 4.280 ;
        RECT 146.930 0.350 147.010 4.280 ;
        RECT 147.850 0.350 147.930 4.280 ;
        RECT 148.770 0.350 148.850 4.280 ;
        RECT 149.690 0.350 149.770 4.280 ;
        RECT 150.610 0.350 150.690 4.280 ;
        RECT 151.530 0.350 151.610 4.280 ;
        RECT 152.450 0.350 152.530 4.280 ;
        RECT 153.370 0.350 153.450 4.280 ;
        RECT 154.290 0.350 154.370 4.280 ;
        RECT 155.210 0.350 155.290 4.280 ;
        RECT 156.130 0.350 156.210 4.280 ;
        RECT 157.050 0.350 157.130 4.280 ;
        RECT 157.970 0.350 158.050 4.280 ;
        RECT 158.890 0.350 158.970 4.280 ;
        RECT 159.810 0.350 159.890 4.280 ;
        RECT 160.730 0.350 160.810 4.280 ;
        RECT 161.650 0.350 161.730 4.280 ;
        RECT 162.570 0.350 162.650 4.280 ;
        RECT 163.490 0.350 163.570 4.280 ;
        RECT 164.410 0.350 164.490 4.280 ;
        RECT 165.330 0.350 165.410 4.280 ;
        RECT 166.250 0.350 166.330 4.280 ;
        RECT 167.170 0.350 167.250 4.280 ;
        RECT 168.090 0.350 168.170 4.280 ;
        RECT 169.010 0.350 169.090 4.280 ;
        RECT 169.930 0.350 170.010 4.280 ;
        RECT 170.850 0.350 170.930 4.280 ;
        RECT 171.770 0.350 171.850 4.280 ;
        RECT 172.690 0.350 172.770 4.280 ;
        RECT 173.610 0.350 173.690 4.280 ;
        RECT 174.530 0.350 174.610 4.280 ;
        RECT 175.450 0.350 175.530 4.280 ;
        RECT 176.370 0.350 176.450 4.280 ;
        RECT 177.290 0.350 177.370 4.280 ;
        RECT 178.210 0.350 178.290 4.280 ;
        RECT 179.130 0.350 179.210 4.280 ;
        RECT 180.050 0.350 180.130 4.280 ;
        RECT 180.970 0.350 181.050 4.280 ;
        RECT 181.890 0.350 181.970 4.280 ;
        RECT 182.810 0.350 182.890 4.280 ;
        RECT 183.730 0.350 183.810 4.280 ;
        RECT 184.650 0.350 184.730 4.280 ;
        RECT 185.570 0.350 185.650 4.280 ;
        RECT 186.490 0.350 186.570 4.280 ;
        RECT 187.410 0.350 187.490 4.280 ;
        RECT 188.330 0.350 188.410 4.280 ;
        RECT 189.250 0.350 189.330 4.280 ;
        RECT 190.170 0.350 190.250 4.280 ;
        RECT 191.090 0.350 191.170 4.280 ;
        RECT 192.010 0.350 192.090 4.280 ;
        RECT 192.930 0.350 193.010 4.280 ;
        RECT 193.850 0.350 193.930 4.280 ;
        RECT 194.770 0.350 194.850 4.280 ;
        RECT 195.690 0.350 195.770 4.280 ;
        RECT 196.610 0.350 196.690 4.280 ;
        RECT 197.530 0.350 197.610 4.280 ;
        RECT 198.450 0.350 198.530 4.280 ;
        RECT 199.370 0.350 199.450 4.280 ;
        RECT 200.290 0.350 200.370 4.280 ;
        RECT 201.210 0.350 201.290 4.280 ;
        RECT 202.130 0.350 202.210 4.280 ;
        RECT 203.050 0.350 203.130 4.280 ;
        RECT 203.970 0.350 204.050 4.280 ;
        RECT 204.890 0.350 204.970 4.280 ;
        RECT 205.810 0.350 205.890 4.280 ;
        RECT 206.730 0.350 206.810 4.280 ;
        RECT 207.650 0.350 207.730 4.280 ;
        RECT 208.570 0.350 208.650 4.280 ;
        RECT 209.490 0.350 209.570 4.280 ;
        RECT 210.410 0.350 210.490 4.280 ;
        RECT 211.330 0.350 211.410 4.280 ;
        RECT 212.250 0.350 212.330 4.280 ;
        RECT 213.170 0.350 213.250 4.280 ;
        RECT 214.090 0.350 214.170 4.280 ;
        RECT 215.010 0.350 215.090 4.280 ;
        RECT 215.930 0.350 216.010 4.280 ;
        RECT 216.850 0.350 216.930 4.280 ;
        RECT 217.770 0.350 217.850 4.280 ;
        RECT 218.690 0.350 218.770 4.280 ;
        RECT 219.610 0.350 219.690 4.280 ;
        RECT 220.530 0.350 220.610 4.280 ;
        RECT 221.450 0.350 221.530 4.280 ;
        RECT 222.370 0.350 222.450 4.280 ;
        RECT 223.290 0.350 223.370 4.280 ;
        RECT 224.210 0.350 224.290 4.280 ;
        RECT 225.130 0.350 225.210 4.280 ;
        RECT 226.050 0.350 226.130 4.280 ;
        RECT 226.970 0.350 227.050 4.280 ;
        RECT 227.890 0.350 227.970 4.280 ;
        RECT 228.810 0.350 228.890 4.280 ;
        RECT 229.730 0.350 229.810 4.280 ;
        RECT 230.650 0.350 230.730 4.280 ;
        RECT 231.570 0.350 231.650 4.280 ;
        RECT 232.490 0.350 232.570 4.280 ;
        RECT 233.410 0.350 233.490 4.280 ;
        RECT 234.330 0.350 234.410 4.280 ;
        RECT 235.250 0.350 235.330 4.280 ;
        RECT 236.170 0.350 236.250 4.280 ;
        RECT 237.090 0.350 237.170 4.280 ;
        RECT 238.010 0.350 238.090 4.280 ;
        RECT 238.930 0.350 239.010 4.280 ;
        RECT 239.850 0.350 239.930 4.280 ;
        RECT 240.770 0.350 240.850 4.280 ;
        RECT 241.690 0.350 241.770 4.280 ;
        RECT 242.610 0.350 242.690 4.280 ;
        RECT 243.530 0.350 243.610 4.280 ;
        RECT 244.450 0.350 244.530 4.280 ;
        RECT 245.370 0.350 245.450 4.280 ;
        RECT 246.290 0.350 246.370 4.280 ;
        RECT 247.210 0.350 247.290 4.280 ;
        RECT 248.130 0.350 248.210 4.280 ;
        RECT 249.050 0.350 249.130 4.280 ;
        RECT 249.970 0.350 250.050 4.280 ;
        RECT 250.890 0.350 250.970 4.280 ;
        RECT 251.810 0.350 251.890 4.280 ;
        RECT 252.730 0.350 252.810 4.280 ;
        RECT 253.650 0.350 253.730 4.280 ;
        RECT 254.570 0.350 254.650 4.280 ;
        RECT 255.490 0.350 255.570 4.280 ;
        RECT 256.410 0.350 256.490 4.280 ;
        RECT 257.330 0.350 257.410 4.280 ;
        RECT 258.250 0.350 258.330 4.280 ;
        RECT 259.170 0.350 259.250 4.280 ;
        RECT 260.090 0.350 260.170 4.280 ;
        RECT 261.010 0.350 261.090 4.280 ;
        RECT 261.930 0.350 262.010 4.280 ;
        RECT 262.850 0.350 262.930 4.280 ;
        RECT 263.770 0.350 263.850 4.280 ;
        RECT 264.690 0.350 264.770 4.280 ;
        RECT 265.610 0.350 265.690 4.280 ;
        RECT 266.530 0.350 266.610 4.280 ;
        RECT 267.450 0.350 267.530 4.280 ;
        RECT 268.370 0.350 268.450 4.280 ;
        RECT 269.290 0.350 269.370 4.280 ;
        RECT 270.210 0.350 270.290 4.280 ;
        RECT 271.130 0.350 271.210 4.280 ;
        RECT 272.050 0.350 272.130 4.280 ;
        RECT 272.970 0.350 273.050 4.280 ;
        RECT 273.890 0.350 273.970 4.280 ;
        RECT 274.810 0.350 274.890 4.280 ;
        RECT 275.730 0.350 275.810 4.280 ;
        RECT 276.650 0.350 276.730 4.280 ;
        RECT 277.570 0.350 277.650 4.280 ;
        RECT 278.490 0.350 278.570 4.280 ;
        RECT 279.410 0.350 279.490 4.280 ;
        RECT 280.330 0.350 280.410 4.280 ;
        RECT 281.250 0.350 281.330 4.280 ;
        RECT 282.170 0.350 282.250 4.280 ;
        RECT 283.090 0.350 283.170 4.280 ;
        RECT 284.010 0.350 284.090 4.280 ;
        RECT 284.930 0.350 285.010 4.280 ;
        RECT 285.850 0.350 285.930 4.280 ;
        RECT 286.770 0.350 286.850 4.280 ;
        RECT 287.690 0.350 287.770 4.280 ;
        RECT 288.610 0.350 288.690 4.280 ;
        RECT 289.530 0.350 289.610 4.280 ;
        RECT 290.450 0.350 290.530 4.280 ;
        RECT 291.370 0.350 291.450 4.280 ;
        RECT 292.290 0.350 292.370 4.280 ;
        RECT 293.210 0.350 293.290 4.280 ;
        RECT 294.130 0.350 294.210 4.280 ;
        RECT 295.050 0.350 295.130 4.280 ;
        RECT 295.970 0.350 296.050 4.280 ;
        RECT 296.890 0.350 296.970 4.280 ;
        RECT 297.810 0.350 297.890 4.280 ;
        RECT 298.730 0.350 298.810 4.280 ;
        RECT 299.650 0.350 299.730 4.280 ;
        RECT 300.570 0.350 300.650 4.280 ;
        RECT 301.490 0.350 301.570 4.280 ;
        RECT 302.410 0.350 302.490 4.280 ;
        RECT 303.330 0.350 303.410 4.280 ;
        RECT 304.250 0.350 304.330 4.280 ;
        RECT 305.170 0.350 305.250 4.280 ;
        RECT 306.090 0.350 306.170 4.280 ;
        RECT 307.010 0.350 307.090 4.280 ;
        RECT 307.930 0.350 308.010 4.280 ;
        RECT 308.850 0.350 308.930 4.280 ;
        RECT 309.770 0.350 309.850 4.280 ;
        RECT 310.690 0.350 310.770 4.280 ;
        RECT 311.610 0.350 311.690 4.280 ;
        RECT 312.530 0.350 312.610 4.280 ;
        RECT 313.450 0.350 313.530 4.280 ;
        RECT 314.370 0.350 314.450 4.280 ;
        RECT 315.290 0.350 315.370 4.280 ;
        RECT 316.210 0.350 316.290 4.280 ;
        RECT 317.130 0.350 317.210 4.280 ;
        RECT 318.050 0.350 318.130 4.280 ;
        RECT 318.970 0.350 319.050 4.280 ;
        RECT 319.890 0.350 319.970 4.280 ;
        RECT 320.810 0.350 320.890 4.280 ;
        RECT 321.730 0.350 321.810 4.280 ;
        RECT 322.650 0.350 322.730 4.280 ;
        RECT 323.570 0.350 323.650 4.280 ;
        RECT 324.490 0.350 324.570 4.280 ;
        RECT 325.410 0.350 325.490 4.280 ;
        RECT 326.330 0.350 326.410 4.280 ;
        RECT 327.250 0.350 327.330 4.280 ;
        RECT 328.170 0.350 328.250 4.280 ;
        RECT 329.090 0.350 329.170 4.280 ;
        RECT 330.010 0.350 330.090 4.280 ;
        RECT 330.930 0.350 331.010 4.280 ;
        RECT 331.850 0.350 331.930 4.280 ;
        RECT 332.770 0.350 332.850 4.280 ;
        RECT 333.690 0.350 333.770 4.280 ;
        RECT 334.610 0.350 334.690 4.280 ;
        RECT 335.530 0.350 335.610 4.280 ;
        RECT 336.450 0.350 336.530 4.280 ;
        RECT 337.370 0.350 337.450 4.280 ;
        RECT 338.290 0.350 338.370 4.280 ;
        RECT 339.210 0.350 339.290 4.280 ;
        RECT 340.130 0.350 340.210 4.280 ;
        RECT 341.050 0.350 341.130 4.280 ;
        RECT 341.970 0.350 342.050 4.280 ;
        RECT 342.890 0.350 342.970 4.280 ;
        RECT 343.810 0.350 343.890 4.280 ;
        RECT 344.730 0.350 344.810 4.280 ;
        RECT 345.650 0.350 345.730 4.280 ;
        RECT 346.570 0.350 346.650 4.280 ;
        RECT 347.490 0.350 347.570 4.280 ;
        RECT 348.410 0.350 348.490 4.280 ;
        RECT 349.330 0.350 349.410 4.280 ;
        RECT 350.250 0.350 350.330 4.280 ;
        RECT 351.170 0.350 351.250 4.280 ;
        RECT 352.090 0.350 352.170 4.280 ;
        RECT 353.010 0.350 353.090 4.280 ;
        RECT 353.930 0.350 354.010 4.280 ;
        RECT 354.850 0.350 354.930 4.280 ;
        RECT 355.770 0.350 355.850 4.280 ;
        RECT 356.690 0.350 356.770 4.280 ;
        RECT 357.610 0.350 357.690 4.280 ;
        RECT 358.530 0.350 358.610 4.280 ;
        RECT 359.450 0.350 359.530 4.280 ;
        RECT 360.370 0.350 360.450 4.280 ;
        RECT 361.290 0.350 361.370 4.280 ;
        RECT 362.210 0.350 362.290 4.280 ;
        RECT 363.130 0.350 363.210 4.280 ;
        RECT 364.050 0.350 364.130 4.280 ;
        RECT 364.970 0.350 365.050 4.280 ;
        RECT 365.890 0.350 365.970 4.280 ;
        RECT 366.810 0.350 366.890 4.280 ;
        RECT 367.730 0.350 367.810 4.280 ;
        RECT 368.650 0.350 368.730 4.280 ;
        RECT 369.570 0.350 369.650 4.280 ;
        RECT 370.490 0.350 370.570 4.280 ;
        RECT 371.410 0.350 371.490 4.280 ;
        RECT 372.330 0.350 372.410 4.280 ;
        RECT 373.250 0.350 373.330 4.280 ;
        RECT 374.170 0.350 374.250 4.280 ;
        RECT 375.090 0.350 375.170 4.280 ;
        RECT 376.010 0.350 376.090 4.280 ;
        RECT 376.930 0.350 377.010 4.280 ;
        RECT 377.850 0.350 377.930 4.280 ;
        RECT 378.770 0.350 378.850 4.280 ;
        RECT 379.690 0.350 379.770 4.280 ;
        RECT 380.610 0.350 380.690 4.280 ;
        RECT 381.530 0.350 381.610 4.280 ;
        RECT 382.450 0.350 382.530 4.280 ;
        RECT 383.370 0.350 383.450 4.280 ;
        RECT 384.290 0.350 384.370 4.280 ;
        RECT 385.210 0.350 385.290 4.280 ;
        RECT 386.130 0.350 386.210 4.280 ;
        RECT 387.050 0.350 387.130 4.280 ;
        RECT 387.970 0.350 388.050 4.280 ;
        RECT 388.890 0.350 388.970 4.280 ;
        RECT 389.810 0.350 389.890 4.280 ;
        RECT 390.730 0.350 390.810 4.280 ;
        RECT 391.650 0.350 391.730 4.280 ;
        RECT 392.570 0.350 392.650 4.280 ;
        RECT 393.490 0.350 393.570 4.280 ;
        RECT 394.410 0.350 394.490 4.280 ;
        RECT 395.330 0.350 395.410 4.280 ;
        RECT 396.250 0.350 396.330 4.280 ;
        RECT 397.170 0.350 397.250 4.280 ;
        RECT 398.090 0.350 398.170 4.280 ;
        RECT 399.010 0.350 399.090 4.280 ;
        RECT 399.930 0.350 400.010 4.280 ;
        RECT 400.850 0.350 400.930 4.280 ;
        RECT 401.770 0.350 401.850 4.280 ;
        RECT 402.690 0.350 402.770 4.280 ;
        RECT 403.610 0.350 403.690 4.280 ;
        RECT 404.530 0.350 404.610 4.280 ;
        RECT 405.450 0.350 405.530 4.280 ;
        RECT 406.370 0.350 406.450 4.280 ;
        RECT 407.290 0.350 407.370 4.280 ;
        RECT 408.210 0.350 408.290 4.280 ;
        RECT 409.130 0.350 409.210 4.280 ;
        RECT 410.050 0.350 410.130 4.280 ;
        RECT 410.970 0.350 411.050 4.280 ;
        RECT 411.890 0.350 411.970 4.280 ;
        RECT 412.810 0.350 412.890 4.280 ;
        RECT 413.730 0.350 413.810 4.280 ;
        RECT 414.650 0.350 414.730 4.280 ;
        RECT 415.570 0.350 450.240 4.280 ;
      LAYER met3 ;
        RECT 12.945 1.535 447.055 454.405 ;
      LAYER met4 ;
        RECT 15.015 10.240 20.640 403.065 ;
        RECT 23.040 10.240 23.940 403.065 ;
        RECT 26.340 10.240 174.240 403.065 ;
        RECT 176.640 10.240 177.540 403.065 ;
        RECT 179.940 10.240 327.840 403.065 ;
        RECT 330.240 10.240 331.140 403.065 ;
        RECT 333.540 10.240 441.305 403.065 ;
        RECT 15.015 1.535 441.305 10.240 ;
  END
END picorv32
END LIBRARY

