VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picorv32
  CLASS BLOCK ;
  FOREIGN picorv32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END clk
  PIN eoi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2448.670 0.000 2448.950 4.000 ;
    END
  END eoi[0]
  PIN eoi[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2536.070 0.000 2536.350 4.000 ;
    END
  END eoi[10]
  PIN eoi[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.810 0.000 2545.090 4.000 ;
    END
  END eoi[11]
  PIN eoi[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.550 0.000 2553.830 4.000 ;
    END
  END eoi[12]
  PIN eoi[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.290 0.000 2562.570 4.000 ;
    END
  END eoi[13]
  PIN eoi[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.030 0.000 2571.310 4.000 ;
    END
  END eoi[14]
  PIN eoi[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.770 0.000 2580.050 4.000 ;
    END
  END eoi[15]
  PIN eoi[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.510 0.000 2588.790 4.000 ;
    END
  END eoi[16]
  PIN eoi[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.250 0.000 2597.530 4.000 ;
    END
  END eoi[17]
  PIN eoi[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.990 0.000 2606.270 4.000 ;
    END
  END eoi[18]
  PIN eoi[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2614.730 0.000 2615.010 4.000 ;
    END
  END eoi[19]
  PIN eoi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2457.410 0.000 2457.690 4.000 ;
    END
  END eoi[1]
  PIN eoi[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2623.470 0.000 2623.750 4.000 ;
    END
  END eoi[20]
  PIN eoi[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.210 0.000 2632.490 4.000 ;
    END
  END eoi[21]
  PIN eoi[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2640.950 0.000 2641.230 4.000 ;
    END
  END eoi[22]
  PIN eoi[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.690 0.000 2649.970 4.000 ;
    END
  END eoi[23]
  PIN eoi[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2658.430 0.000 2658.710 4.000 ;
    END
  END eoi[24]
  PIN eoi[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.170 0.000 2667.450 4.000 ;
    END
  END eoi[25]
  PIN eoi[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.910 0.000 2676.190 4.000 ;
    END
  END eoi[26]
  PIN eoi[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.650 0.000 2684.930 4.000 ;
    END
  END eoi[27]
  PIN eoi[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.390 0.000 2693.670 4.000 ;
    END
  END eoi[28]
  PIN eoi[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.130 0.000 2702.410 4.000 ;
    END
  END eoi[29]
  PIN eoi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.150 0.000 2466.430 4.000 ;
    END
  END eoi[2]
  PIN eoi[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2710.870 0.000 2711.150 4.000 ;
    END
  END eoi[30]
  PIN eoi[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2719.610 0.000 2719.890 4.000 ;
    END
  END eoi[31]
  PIN eoi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2474.890 0.000 2475.170 4.000 ;
    END
  END eoi[3]
  PIN eoi[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.630 0.000 2483.910 4.000 ;
    END
  END eoi[4]
  PIN eoi[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.370 0.000 2492.650 4.000 ;
    END
  END eoi[5]
  PIN eoi[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2501.110 0.000 2501.390 4.000 ;
    END
  END eoi[6]
  PIN eoi[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2509.850 0.000 2510.130 4.000 ;
    END
  END eoi[7]
  PIN eoi[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.590 0.000 2518.870 4.000 ;
    END
  END eoi[8]
  PIN eoi[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.330 0.000 2527.610 4.000 ;
    END
  END eoi[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END irq[15]
  PIN irq[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END irq[16]
  PIN irq[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END irq[17]
  PIN irq[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END irq[18]
  PIN irq[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END irq[19]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END irq[1]
  PIN irq[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END irq[20]
  PIN irq[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END irq[21]
  PIN irq[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END irq[22]
  PIN irq[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END irq[23]
  PIN irq[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END irq[24]
  PIN irq[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END irq[25]
  PIN irq[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END irq[26]
  PIN irq[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END irq[27]
  PIN irq[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END irq[28]
  PIN irq[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END irq[29]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END irq[2]
  PIN irq[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END irq[30]
  PIN irq[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END irq[31]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END irq[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.920 4.000 1745.520 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1486.520 4.000 1487.120 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.680 4.000 1461.280 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.160 4.000 1383.760 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1357.320 4.000 1357.920 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.800 4.000 1280.400 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.960 4.000 1254.560 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 4.000 1719.680 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.120 4.000 1228.720 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 4.000 1202.880 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1150.600 4.000 1151.200 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.080 4.000 1073.680 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 995.560 4.000 996.160 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1667.400 4.000 1668.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1641.560 4.000 1642.160 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1615.720 4.000 1616.320 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.880 4.000 1590.480 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1538.200 4.000 1538.800 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1512.360 4.000 1512.960 ;
    END
  END mem_addr[9]
  PIN mem_instr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2728.350 0.000 2728.630 4.000 ;
    END
  END mem_instr
  PIN mem_la_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.970 0.000 1531.250 4.000 ;
    END
  END mem_la_addr[0]
  PIN mem_la_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1740.730 0.000 1741.010 4.000 ;
    END
  END mem_la_addr[10]
  PIN mem_la_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END mem_la_addr[11]
  PIN mem_la_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1775.690 0.000 1775.970 4.000 ;
    END
  END mem_la_addr[12]
  PIN mem_la_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1793.170 0.000 1793.450 4.000 ;
    END
  END mem_la_addr[13]
  PIN mem_la_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1810.650 0.000 1810.930 4.000 ;
    END
  END mem_la_addr[14]
  PIN mem_la_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1828.130 0.000 1828.410 4.000 ;
    END
  END mem_la_addr[15]
  PIN mem_la_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1845.610 0.000 1845.890 4.000 ;
    END
  END mem_la_addr[16]
  PIN mem_la_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1863.090 0.000 1863.370 4.000 ;
    END
  END mem_la_addr[17]
  PIN mem_la_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END mem_la_addr[18]
  PIN mem_la_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1898.050 0.000 1898.330 4.000 ;
    END
  END mem_la_addr[19]
  PIN mem_la_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 0.000 1557.470 4.000 ;
    END
  END mem_la_addr[1]
  PIN mem_la_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END mem_la_addr[20]
  PIN mem_la_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1933.010 0.000 1933.290 4.000 ;
    END
  END mem_la_addr[21]
  PIN mem_la_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1950.490 0.000 1950.770 4.000 ;
    END
  END mem_la_addr[22]
  PIN mem_la_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1967.970 0.000 1968.250 4.000 ;
    END
  END mem_la_addr[23]
  PIN mem_la_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1985.450 0.000 1985.730 4.000 ;
    END
  END mem_la_addr[24]
  PIN mem_la_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2002.930 0.000 2003.210 4.000 ;
    END
  END mem_la_addr[25]
  PIN mem_la_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2020.410 0.000 2020.690 4.000 ;
    END
  END mem_la_addr[26]
  PIN mem_la_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2037.890 0.000 2038.170 4.000 ;
    END
  END mem_la_addr[27]
  PIN mem_la_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2055.370 0.000 2055.650 4.000 ;
    END
  END mem_la_addr[28]
  PIN mem_la_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2072.850 0.000 2073.130 4.000 ;
    END
  END mem_la_addr[29]
  PIN mem_la_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1583.410 0.000 1583.690 4.000 ;
    END
  END mem_la_addr[2]
  PIN mem_la_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2090.330 0.000 2090.610 4.000 ;
    END
  END mem_la_addr[30]
  PIN mem_la_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2107.810 0.000 2108.090 4.000 ;
    END
  END mem_la_addr[31]
  PIN mem_la_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1609.630 0.000 1609.910 4.000 ;
    END
  END mem_la_addr[3]
  PIN mem_la_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END mem_la_addr[4]
  PIN mem_la_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1653.330 0.000 1653.610 4.000 ;
    END
  END mem_la_addr[5]
  PIN mem_la_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END mem_la_addr[6]
  PIN mem_la_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1688.290 0.000 1688.570 4.000 ;
    END
  END mem_la_addr[7]
  PIN mem_la_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1705.770 0.000 1706.050 4.000 ;
    END
  END mem_la_addr[8]
  PIN mem_la_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1723.250 0.000 1723.530 4.000 ;
    END
  END mem_la_addr[9]
  PIN mem_la_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END mem_la_read
  PIN mem_la_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END mem_la_wdata[0]
  PIN mem_la_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 4.000 ;
    END
  END mem_la_wdata[10]
  PIN mem_la_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1766.950 0.000 1767.230 4.000 ;
    END
  END mem_la_wdata[11]
  PIN mem_la_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1784.430 0.000 1784.710 4.000 ;
    END
  END mem_la_wdata[12]
  PIN mem_la_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 4.000 ;
    END
  END mem_la_wdata[13]
  PIN mem_la_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1819.390 0.000 1819.670 4.000 ;
    END
  END mem_la_wdata[14]
  PIN mem_la_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1836.870 0.000 1837.150 4.000 ;
    END
  END mem_la_wdata[15]
  PIN mem_la_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1854.350 0.000 1854.630 4.000 ;
    END
  END mem_la_wdata[16]
  PIN mem_la_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1871.830 0.000 1872.110 4.000 ;
    END
  END mem_la_wdata[17]
  PIN mem_la_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1889.310 0.000 1889.590 4.000 ;
    END
  END mem_la_wdata[18]
  PIN mem_la_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1906.790 0.000 1907.070 4.000 ;
    END
  END mem_la_wdata[19]
  PIN mem_la_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1565.930 0.000 1566.210 4.000 ;
    END
  END mem_la_wdata[1]
  PIN mem_la_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1924.270 0.000 1924.550 4.000 ;
    END
  END mem_la_wdata[20]
  PIN mem_la_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1941.750 0.000 1942.030 4.000 ;
    END
  END mem_la_wdata[21]
  PIN mem_la_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END mem_la_wdata[22]
  PIN mem_la_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1976.710 0.000 1976.990 4.000 ;
    END
  END mem_la_wdata[23]
  PIN mem_la_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1994.190 0.000 1994.470 4.000 ;
    END
  END mem_la_wdata[24]
  PIN mem_la_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2011.670 0.000 2011.950 4.000 ;
    END
  END mem_la_wdata[25]
  PIN mem_la_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2029.150 0.000 2029.430 4.000 ;
    END
  END mem_la_wdata[26]
  PIN mem_la_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2046.630 0.000 2046.910 4.000 ;
    END
  END mem_la_wdata[27]
  PIN mem_la_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END mem_la_wdata[28]
  PIN mem_la_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2081.590 0.000 2081.870 4.000 ;
    END
  END mem_la_wdata[29]
  PIN mem_la_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1592.150 0.000 1592.430 4.000 ;
    END
  END mem_la_wdata[2]
  PIN mem_la_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2099.070 0.000 2099.350 4.000 ;
    END
  END mem_la_wdata[30]
  PIN mem_la_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2116.550 0.000 2116.830 4.000 ;
    END
  END mem_la_wdata[31]
  PIN mem_la_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1618.370 0.000 1618.650 4.000 ;
    END
  END mem_la_wdata[3]
  PIN mem_la_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1644.590 0.000 1644.870 4.000 ;
    END
  END mem_la_wdata[4]
  PIN mem_la_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1662.070 0.000 1662.350 4.000 ;
    END
  END mem_la_wdata[5]
  PIN mem_la_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1679.550 0.000 1679.830 4.000 ;
    END
  END mem_la_wdata[6]
  PIN mem_la_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END mem_la_wdata[7]
  PIN mem_la_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1714.510 0.000 1714.790 4.000 ;
    END
  END mem_la_wdata[8]
  PIN mem_la_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1731.990 0.000 1732.270 4.000 ;
    END
  END mem_la_wdata[9]
  PIN mem_la_write
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1522.230 0.000 1522.510 4.000 ;
    END
  END mem_la_write
  PIN mem_la_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1548.450 0.000 1548.730 4.000 ;
    END
  END mem_la_wstrb[0]
  PIN mem_la_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END mem_la_wstrb[1]
  PIN mem_la_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END mem_la_wstrb[2]
  PIN mem_la_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1627.110 0.000 1627.390 4.000 ;
    END
  END mem_la_wstrb[3]
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 35.400 2800.000 36.000 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 579.400 2800.000 580.000 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 633.800 2800.000 634.400 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 688.200 2800.000 688.800 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 742.600 2800.000 743.200 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 797.000 2800.000 797.600 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 851.400 2800.000 852.000 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 905.800 2800.000 906.400 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 960.200 2800.000 960.800 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1014.600 2800.000 1015.200 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1069.000 2800.000 1069.600 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 89.800 2800.000 90.400 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1123.400 2800.000 1124.000 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1177.800 2800.000 1178.400 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1232.200 2800.000 1232.800 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1286.600 2800.000 1287.200 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1341.000 2800.000 1341.600 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1395.400 2800.000 1396.000 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1449.800 2800.000 1450.400 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1504.200 2800.000 1504.800 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1558.600 2800.000 1559.200 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1613.000 2800.000 1613.600 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 144.200 2800.000 144.800 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1667.400 2800.000 1668.000 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1721.800 2800.000 1722.400 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 198.600 2800.000 199.200 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 253.000 2800.000 253.600 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 307.400 2800.000 308.000 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 361.800 2800.000 362.400 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 416.200 2800.000 416.800 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 470.600 2800.000 471.200 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 525.000 2800.000 525.600 ;
    END
  END mem_rdata[9]
  PIN mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 2737.090 0.000 2737.370 4.000 ;
    END
  END mem_ready
  PIN mem_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2745.830 0.000 2746.110 4.000 ;
    END
  END mem_valid
  PIN mem_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END mem_wdata[9]
  PIN mem_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END mem_wstrb[0]
  PIN mem_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mem_wstrb[1]
  PIN mem_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END mem_wstrb[2]
  PIN mem_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mem_wstrb[3]
  PIN pcpi_insn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 0.000 989.370 4.000 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 0.000 1199.130 4.000 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 0.000 1234.090 4.000 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 0.000 1304.010 4.000 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.690 0.000 1338.970 4.000 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 0.000 1373.930 4.000 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 0.000 1443.850 4.000 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.790 0.000 1033.070 4.000 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 0.000 1172.910 4.000 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 0.000 1242.830 4.000 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 0.000 1312.750 4.000 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.430 0.000 1347.710 4.000 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 0.000 1382.670 4.000 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 0.000 1417.630 4.000 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.270 0.000 1487.550 4.000 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 0.000 648.510 4.000 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1041.530 0.000 1041.810 4.000 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1111.450 0.000 1111.730 4.000 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1181.370 0.000 1181.650 4.000 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1251.290 0.000 1251.570 4.000 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1286.250 0.000 1286.530 4.000 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1321.210 0.000 1321.490 4.000 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1356.170 0.000 1356.450 4.000 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 4.000 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1496.010 0.000 1496.290 4.000 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 875.470 0.000 875.750 4.000 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1225.070 0.000 1225.350 4.000 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 4.000 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1364.910 0.000 1365.190 4.000 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1434.830 0.000 1435.110 4.000 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1469.790 0.000 1470.070 4.000 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1504.750 0.000 1505.030 4.000 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END resetn
  PIN trace_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.030 0.000 2134.310 4.000 ;
    END
  END trace_data[0]
  PIN trace_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.430 0.000 2221.710 4.000 ;
    END
  END trace_data[10]
  PIN trace_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.170 0.000 2230.450 4.000 ;
    END
  END trace_data[11]
  PIN trace_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.910 0.000 2239.190 4.000 ;
    END
  END trace_data[12]
  PIN trace_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END trace_data[13]
  PIN trace_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.390 0.000 2256.670 4.000 ;
    END
  END trace_data[14]
  PIN trace_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2265.130 0.000 2265.410 4.000 ;
    END
  END trace_data[15]
  PIN trace_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.870 0.000 2274.150 4.000 ;
    END
  END trace_data[16]
  PIN trace_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.610 0.000 2282.890 4.000 ;
    END
  END trace_data[17]
  PIN trace_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2291.350 0.000 2291.630 4.000 ;
    END
  END trace_data[18]
  PIN trace_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2300.090 0.000 2300.370 4.000 ;
    END
  END trace_data[19]
  PIN trace_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.770 0.000 2143.050 4.000 ;
    END
  END trace_data[1]
  PIN trace_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.830 0.000 2309.110 4.000 ;
    END
  END trace_data[20]
  PIN trace_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.570 0.000 2317.850 4.000 ;
    END
  END trace_data[21]
  PIN trace_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2326.310 0.000 2326.590 4.000 ;
    END
  END trace_data[22]
  PIN trace_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.050 0.000 2335.330 4.000 ;
    END
  END trace_data[23]
  PIN trace_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.790 0.000 2344.070 4.000 ;
    END
  END trace_data[24]
  PIN trace_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.530 0.000 2352.810 4.000 ;
    END
  END trace_data[25]
  PIN trace_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.270 0.000 2361.550 4.000 ;
    END
  END trace_data[26]
  PIN trace_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 0.000 2370.290 4.000 ;
    END
  END trace_data[27]
  PIN trace_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.750 0.000 2379.030 4.000 ;
    END
  END trace_data[28]
  PIN trace_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.490 0.000 2387.770 4.000 ;
    END
  END trace_data[29]
  PIN trace_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.510 0.000 2151.790 4.000 ;
    END
  END trace_data[2]
  PIN trace_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.230 0.000 2396.510 4.000 ;
    END
  END trace_data[30]
  PIN trace_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.970 0.000 2405.250 4.000 ;
    END
  END trace_data[31]
  PIN trace_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 4.000 ;
    END
  END trace_data[32]
  PIN trace_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.450 0.000 2422.730 4.000 ;
    END
  END trace_data[33]
  PIN trace_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 4.000 ;
    END
  END trace_data[34]
  PIN trace_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.930 0.000 2440.210 4.000 ;
    END
  END trace_data[35]
  PIN trace_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.250 0.000 2160.530 4.000 ;
    END
  END trace_data[3]
  PIN trace_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 4.000 ;
    END
  END trace_data[4]
  PIN trace_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.730 0.000 2178.010 4.000 ;
    END
  END trace_data[5]
  PIN trace_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 0.000 2186.750 4.000 ;
    END
  END trace_data[6]
  PIN trace_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.210 0.000 2195.490 4.000 ;
    END
  END trace_data[7]
  PIN trace_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.950 0.000 2204.230 4.000 ;
    END
  END trace_data[8]
  PIN trace_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.690 0.000 2212.970 4.000 ;
    END
  END trace_data[9]
  PIN trace_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 4.000 ;
    END
  END trace_valid
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END trap
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 1.400 2794.340 1749.200 ;
      LAYER met2 ;
        RECT 4.690 4.280 2792.560 1749.145 ;
        RECT 4.690 1.370 53.630 4.280 ;
        RECT 54.470 1.370 62.370 4.280 ;
        RECT 63.210 1.370 71.110 4.280 ;
        RECT 71.950 1.370 79.850 4.280 ;
        RECT 80.690 1.370 88.590 4.280 ;
        RECT 89.430 1.370 97.330 4.280 ;
        RECT 98.170 1.370 106.070 4.280 ;
        RECT 106.910 1.370 114.810 4.280 ;
        RECT 115.650 1.370 123.550 4.280 ;
        RECT 124.390 1.370 132.290 4.280 ;
        RECT 133.130 1.370 141.030 4.280 ;
        RECT 141.870 1.370 149.770 4.280 ;
        RECT 150.610 1.370 158.510 4.280 ;
        RECT 159.350 1.370 167.250 4.280 ;
        RECT 168.090 1.370 175.990 4.280 ;
        RECT 176.830 1.370 184.730 4.280 ;
        RECT 185.570 1.370 193.470 4.280 ;
        RECT 194.310 1.370 202.210 4.280 ;
        RECT 203.050 1.370 210.950 4.280 ;
        RECT 211.790 1.370 219.690 4.280 ;
        RECT 220.530 1.370 228.430 4.280 ;
        RECT 229.270 1.370 237.170 4.280 ;
        RECT 238.010 1.370 245.910 4.280 ;
        RECT 246.750 1.370 254.650 4.280 ;
        RECT 255.490 1.370 263.390 4.280 ;
        RECT 264.230 1.370 272.130 4.280 ;
        RECT 272.970 1.370 280.870 4.280 ;
        RECT 281.710 1.370 289.610 4.280 ;
        RECT 290.450 1.370 298.350 4.280 ;
        RECT 299.190 1.370 307.090 4.280 ;
        RECT 307.930 1.370 315.830 4.280 ;
        RECT 316.670 1.370 324.570 4.280 ;
        RECT 325.410 1.370 333.310 4.280 ;
        RECT 334.150 1.370 342.050 4.280 ;
        RECT 342.890 1.370 350.790 4.280 ;
        RECT 351.630 1.370 359.530 4.280 ;
        RECT 360.370 1.370 368.270 4.280 ;
        RECT 369.110 1.370 377.010 4.280 ;
        RECT 377.850 1.370 385.750 4.280 ;
        RECT 386.590 1.370 394.490 4.280 ;
        RECT 395.330 1.370 403.230 4.280 ;
        RECT 404.070 1.370 411.970 4.280 ;
        RECT 412.810 1.370 420.710 4.280 ;
        RECT 421.550 1.370 429.450 4.280 ;
        RECT 430.290 1.370 438.190 4.280 ;
        RECT 439.030 1.370 446.930 4.280 ;
        RECT 447.770 1.370 455.670 4.280 ;
        RECT 456.510 1.370 464.410 4.280 ;
        RECT 465.250 1.370 473.150 4.280 ;
        RECT 473.990 1.370 481.890 4.280 ;
        RECT 482.730 1.370 490.630 4.280 ;
        RECT 491.470 1.370 499.370 4.280 ;
        RECT 500.210 1.370 508.110 4.280 ;
        RECT 508.950 1.370 516.850 4.280 ;
        RECT 517.690 1.370 525.590 4.280 ;
        RECT 526.430 1.370 534.330 4.280 ;
        RECT 535.170 1.370 543.070 4.280 ;
        RECT 543.910 1.370 551.810 4.280 ;
        RECT 552.650 1.370 560.550 4.280 ;
        RECT 561.390 1.370 569.290 4.280 ;
        RECT 570.130 1.370 578.030 4.280 ;
        RECT 578.870 1.370 586.770 4.280 ;
        RECT 587.610 1.370 595.510 4.280 ;
        RECT 596.350 1.370 604.250 4.280 ;
        RECT 605.090 1.370 612.990 4.280 ;
        RECT 613.830 1.370 621.730 4.280 ;
        RECT 622.570 1.370 630.470 4.280 ;
        RECT 631.310 1.370 639.210 4.280 ;
        RECT 640.050 1.370 647.950 4.280 ;
        RECT 648.790 1.370 656.690 4.280 ;
        RECT 657.530 1.370 665.430 4.280 ;
        RECT 666.270 1.370 674.170 4.280 ;
        RECT 675.010 1.370 682.910 4.280 ;
        RECT 683.750 1.370 691.650 4.280 ;
        RECT 692.490 1.370 700.390 4.280 ;
        RECT 701.230 1.370 709.130 4.280 ;
        RECT 709.970 1.370 717.870 4.280 ;
        RECT 718.710 1.370 726.610 4.280 ;
        RECT 727.450 1.370 735.350 4.280 ;
        RECT 736.190 1.370 744.090 4.280 ;
        RECT 744.930 1.370 752.830 4.280 ;
        RECT 753.670 1.370 761.570 4.280 ;
        RECT 762.410 1.370 770.310 4.280 ;
        RECT 771.150 1.370 779.050 4.280 ;
        RECT 779.890 1.370 787.790 4.280 ;
        RECT 788.630 1.370 796.530 4.280 ;
        RECT 797.370 1.370 805.270 4.280 ;
        RECT 806.110 1.370 814.010 4.280 ;
        RECT 814.850 1.370 822.750 4.280 ;
        RECT 823.590 1.370 831.490 4.280 ;
        RECT 832.330 1.370 840.230 4.280 ;
        RECT 841.070 1.370 848.970 4.280 ;
        RECT 849.810 1.370 857.710 4.280 ;
        RECT 858.550 1.370 866.450 4.280 ;
        RECT 867.290 1.370 875.190 4.280 ;
        RECT 876.030 1.370 883.930 4.280 ;
        RECT 884.770 1.370 892.670 4.280 ;
        RECT 893.510 1.370 901.410 4.280 ;
        RECT 902.250 1.370 910.150 4.280 ;
        RECT 910.990 1.370 918.890 4.280 ;
        RECT 919.730 1.370 927.630 4.280 ;
        RECT 928.470 1.370 936.370 4.280 ;
        RECT 937.210 1.370 945.110 4.280 ;
        RECT 945.950 1.370 953.850 4.280 ;
        RECT 954.690 1.370 962.590 4.280 ;
        RECT 963.430 1.370 971.330 4.280 ;
        RECT 972.170 1.370 980.070 4.280 ;
        RECT 980.910 1.370 988.810 4.280 ;
        RECT 989.650 1.370 997.550 4.280 ;
        RECT 998.390 1.370 1006.290 4.280 ;
        RECT 1007.130 1.370 1015.030 4.280 ;
        RECT 1015.870 1.370 1023.770 4.280 ;
        RECT 1024.610 1.370 1032.510 4.280 ;
        RECT 1033.350 1.370 1041.250 4.280 ;
        RECT 1042.090 1.370 1049.990 4.280 ;
        RECT 1050.830 1.370 1058.730 4.280 ;
        RECT 1059.570 1.370 1067.470 4.280 ;
        RECT 1068.310 1.370 1076.210 4.280 ;
        RECT 1077.050 1.370 1084.950 4.280 ;
        RECT 1085.790 1.370 1093.690 4.280 ;
        RECT 1094.530 1.370 1102.430 4.280 ;
        RECT 1103.270 1.370 1111.170 4.280 ;
        RECT 1112.010 1.370 1119.910 4.280 ;
        RECT 1120.750 1.370 1128.650 4.280 ;
        RECT 1129.490 1.370 1137.390 4.280 ;
        RECT 1138.230 1.370 1146.130 4.280 ;
        RECT 1146.970 1.370 1154.870 4.280 ;
        RECT 1155.710 1.370 1163.610 4.280 ;
        RECT 1164.450 1.370 1172.350 4.280 ;
        RECT 1173.190 1.370 1181.090 4.280 ;
        RECT 1181.930 1.370 1189.830 4.280 ;
        RECT 1190.670 1.370 1198.570 4.280 ;
        RECT 1199.410 1.370 1207.310 4.280 ;
        RECT 1208.150 1.370 1216.050 4.280 ;
        RECT 1216.890 1.370 1224.790 4.280 ;
        RECT 1225.630 1.370 1233.530 4.280 ;
        RECT 1234.370 1.370 1242.270 4.280 ;
        RECT 1243.110 1.370 1251.010 4.280 ;
        RECT 1251.850 1.370 1259.750 4.280 ;
        RECT 1260.590 1.370 1268.490 4.280 ;
        RECT 1269.330 1.370 1277.230 4.280 ;
        RECT 1278.070 1.370 1285.970 4.280 ;
        RECT 1286.810 1.370 1294.710 4.280 ;
        RECT 1295.550 1.370 1303.450 4.280 ;
        RECT 1304.290 1.370 1312.190 4.280 ;
        RECT 1313.030 1.370 1320.930 4.280 ;
        RECT 1321.770 1.370 1329.670 4.280 ;
        RECT 1330.510 1.370 1338.410 4.280 ;
        RECT 1339.250 1.370 1347.150 4.280 ;
        RECT 1347.990 1.370 1355.890 4.280 ;
        RECT 1356.730 1.370 1364.630 4.280 ;
        RECT 1365.470 1.370 1373.370 4.280 ;
        RECT 1374.210 1.370 1382.110 4.280 ;
        RECT 1382.950 1.370 1390.850 4.280 ;
        RECT 1391.690 1.370 1399.590 4.280 ;
        RECT 1400.430 1.370 1408.330 4.280 ;
        RECT 1409.170 1.370 1417.070 4.280 ;
        RECT 1417.910 1.370 1425.810 4.280 ;
        RECT 1426.650 1.370 1434.550 4.280 ;
        RECT 1435.390 1.370 1443.290 4.280 ;
        RECT 1444.130 1.370 1452.030 4.280 ;
        RECT 1452.870 1.370 1460.770 4.280 ;
        RECT 1461.610 1.370 1469.510 4.280 ;
        RECT 1470.350 1.370 1478.250 4.280 ;
        RECT 1479.090 1.370 1486.990 4.280 ;
        RECT 1487.830 1.370 1495.730 4.280 ;
        RECT 1496.570 1.370 1504.470 4.280 ;
        RECT 1505.310 1.370 1513.210 4.280 ;
        RECT 1514.050 1.370 1521.950 4.280 ;
        RECT 1522.790 1.370 1530.690 4.280 ;
        RECT 1531.530 1.370 1539.430 4.280 ;
        RECT 1540.270 1.370 1548.170 4.280 ;
        RECT 1549.010 1.370 1556.910 4.280 ;
        RECT 1557.750 1.370 1565.650 4.280 ;
        RECT 1566.490 1.370 1574.390 4.280 ;
        RECT 1575.230 1.370 1583.130 4.280 ;
        RECT 1583.970 1.370 1591.870 4.280 ;
        RECT 1592.710 1.370 1600.610 4.280 ;
        RECT 1601.450 1.370 1609.350 4.280 ;
        RECT 1610.190 1.370 1618.090 4.280 ;
        RECT 1618.930 1.370 1626.830 4.280 ;
        RECT 1627.670 1.370 1635.570 4.280 ;
        RECT 1636.410 1.370 1644.310 4.280 ;
        RECT 1645.150 1.370 1653.050 4.280 ;
        RECT 1653.890 1.370 1661.790 4.280 ;
        RECT 1662.630 1.370 1670.530 4.280 ;
        RECT 1671.370 1.370 1679.270 4.280 ;
        RECT 1680.110 1.370 1688.010 4.280 ;
        RECT 1688.850 1.370 1696.750 4.280 ;
        RECT 1697.590 1.370 1705.490 4.280 ;
        RECT 1706.330 1.370 1714.230 4.280 ;
        RECT 1715.070 1.370 1722.970 4.280 ;
        RECT 1723.810 1.370 1731.710 4.280 ;
        RECT 1732.550 1.370 1740.450 4.280 ;
        RECT 1741.290 1.370 1749.190 4.280 ;
        RECT 1750.030 1.370 1757.930 4.280 ;
        RECT 1758.770 1.370 1766.670 4.280 ;
        RECT 1767.510 1.370 1775.410 4.280 ;
        RECT 1776.250 1.370 1784.150 4.280 ;
        RECT 1784.990 1.370 1792.890 4.280 ;
        RECT 1793.730 1.370 1801.630 4.280 ;
        RECT 1802.470 1.370 1810.370 4.280 ;
        RECT 1811.210 1.370 1819.110 4.280 ;
        RECT 1819.950 1.370 1827.850 4.280 ;
        RECT 1828.690 1.370 1836.590 4.280 ;
        RECT 1837.430 1.370 1845.330 4.280 ;
        RECT 1846.170 1.370 1854.070 4.280 ;
        RECT 1854.910 1.370 1862.810 4.280 ;
        RECT 1863.650 1.370 1871.550 4.280 ;
        RECT 1872.390 1.370 1880.290 4.280 ;
        RECT 1881.130 1.370 1889.030 4.280 ;
        RECT 1889.870 1.370 1897.770 4.280 ;
        RECT 1898.610 1.370 1906.510 4.280 ;
        RECT 1907.350 1.370 1915.250 4.280 ;
        RECT 1916.090 1.370 1923.990 4.280 ;
        RECT 1924.830 1.370 1932.730 4.280 ;
        RECT 1933.570 1.370 1941.470 4.280 ;
        RECT 1942.310 1.370 1950.210 4.280 ;
        RECT 1951.050 1.370 1958.950 4.280 ;
        RECT 1959.790 1.370 1967.690 4.280 ;
        RECT 1968.530 1.370 1976.430 4.280 ;
        RECT 1977.270 1.370 1985.170 4.280 ;
        RECT 1986.010 1.370 1993.910 4.280 ;
        RECT 1994.750 1.370 2002.650 4.280 ;
        RECT 2003.490 1.370 2011.390 4.280 ;
        RECT 2012.230 1.370 2020.130 4.280 ;
        RECT 2020.970 1.370 2028.870 4.280 ;
        RECT 2029.710 1.370 2037.610 4.280 ;
        RECT 2038.450 1.370 2046.350 4.280 ;
        RECT 2047.190 1.370 2055.090 4.280 ;
        RECT 2055.930 1.370 2063.830 4.280 ;
        RECT 2064.670 1.370 2072.570 4.280 ;
        RECT 2073.410 1.370 2081.310 4.280 ;
        RECT 2082.150 1.370 2090.050 4.280 ;
        RECT 2090.890 1.370 2098.790 4.280 ;
        RECT 2099.630 1.370 2107.530 4.280 ;
        RECT 2108.370 1.370 2116.270 4.280 ;
        RECT 2117.110 1.370 2125.010 4.280 ;
        RECT 2125.850 1.370 2133.750 4.280 ;
        RECT 2134.590 1.370 2142.490 4.280 ;
        RECT 2143.330 1.370 2151.230 4.280 ;
        RECT 2152.070 1.370 2159.970 4.280 ;
        RECT 2160.810 1.370 2168.710 4.280 ;
        RECT 2169.550 1.370 2177.450 4.280 ;
        RECT 2178.290 1.370 2186.190 4.280 ;
        RECT 2187.030 1.370 2194.930 4.280 ;
        RECT 2195.770 1.370 2203.670 4.280 ;
        RECT 2204.510 1.370 2212.410 4.280 ;
        RECT 2213.250 1.370 2221.150 4.280 ;
        RECT 2221.990 1.370 2229.890 4.280 ;
        RECT 2230.730 1.370 2238.630 4.280 ;
        RECT 2239.470 1.370 2247.370 4.280 ;
        RECT 2248.210 1.370 2256.110 4.280 ;
        RECT 2256.950 1.370 2264.850 4.280 ;
        RECT 2265.690 1.370 2273.590 4.280 ;
        RECT 2274.430 1.370 2282.330 4.280 ;
        RECT 2283.170 1.370 2291.070 4.280 ;
        RECT 2291.910 1.370 2299.810 4.280 ;
        RECT 2300.650 1.370 2308.550 4.280 ;
        RECT 2309.390 1.370 2317.290 4.280 ;
        RECT 2318.130 1.370 2326.030 4.280 ;
        RECT 2326.870 1.370 2334.770 4.280 ;
        RECT 2335.610 1.370 2343.510 4.280 ;
        RECT 2344.350 1.370 2352.250 4.280 ;
        RECT 2353.090 1.370 2360.990 4.280 ;
        RECT 2361.830 1.370 2369.730 4.280 ;
        RECT 2370.570 1.370 2378.470 4.280 ;
        RECT 2379.310 1.370 2387.210 4.280 ;
        RECT 2388.050 1.370 2395.950 4.280 ;
        RECT 2396.790 1.370 2404.690 4.280 ;
        RECT 2405.530 1.370 2413.430 4.280 ;
        RECT 2414.270 1.370 2422.170 4.280 ;
        RECT 2423.010 1.370 2430.910 4.280 ;
        RECT 2431.750 1.370 2439.650 4.280 ;
        RECT 2440.490 1.370 2448.390 4.280 ;
        RECT 2449.230 1.370 2457.130 4.280 ;
        RECT 2457.970 1.370 2465.870 4.280 ;
        RECT 2466.710 1.370 2474.610 4.280 ;
        RECT 2475.450 1.370 2483.350 4.280 ;
        RECT 2484.190 1.370 2492.090 4.280 ;
        RECT 2492.930 1.370 2500.830 4.280 ;
        RECT 2501.670 1.370 2509.570 4.280 ;
        RECT 2510.410 1.370 2518.310 4.280 ;
        RECT 2519.150 1.370 2527.050 4.280 ;
        RECT 2527.890 1.370 2535.790 4.280 ;
        RECT 2536.630 1.370 2544.530 4.280 ;
        RECT 2545.370 1.370 2553.270 4.280 ;
        RECT 2554.110 1.370 2562.010 4.280 ;
        RECT 2562.850 1.370 2570.750 4.280 ;
        RECT 2571.590 1.370 2579.490 4.280 ;
        RECT 2580.330 1.370 2588.230 4.280 ;
        RECT 2589.070 1.370 2596.970 4.280 ;
        RECT 2597.810 1.370 2605.710 4.280 ;
        RECT 2606.550 1.370 2614.450 4.280 ;
        RECT 2615.290 1.370 2623.190 4.280 ;
        RECT 2624.030 1.370 2631.930 4.280 ;
        RECT 2632.770 1.370 2640.670 4.280 ;
        RECT 2641.510 1.370 2649.410 4.280 ;
        RECT 2650.250 1.370 2658.150 4.280 ;
        RECT 2658.990 1.370 2666.890 4.280 ;
        RECT 2667.730 1.370 2675.630 4.280 ;
        RECT 2676.470 1.370 2684.370 4.280 ;
        RECT 2685.210 1.370 2693.110 4.280 ;
        RECT 2693.950 1.370 2701.850 4.280 ;
        RECT 2702.690 1.370 2710.590 4.280 ;
        RECT 2711.430 1.370 2719.330 4.280 ;
        RECT 2720.170 1.370 2728.070 4.280 ;
        RECT 2728.910 1.370 2736.810 4.280 ;
        RECT 2737.650 1.370 2745.550 4.280 ;
        RECT 2746.390 1.370 2792.560 4.280 ;
      LAYER met3 ;
        RECT 4.000 1745.920 2796.000 1749.125 ;
        RECT 4.400 1744.520 2796.000 1745.920 ;
        RECT 4.000 1722.800 2796.000 1744.520 ;
        RECT 4.000 1721.400 2795.600 1722.800 ;
        RECT 4.000 1720.080 2796.000 1721.400 ;
        RECT 4.400 1718.680 2796.000 1720.080 ;
        RECT 4.000 1694.240 2796.000 1718.680 ;
        RECT 4.400 1692.840 2796.000 1694.240 ;
        RECT 4.000 1668.400 2796.000 1692.840 ;
        RECT 4.400 1667.000 2795.600 1668.400 ;
        RECT 4.000 1642.560 2796.000 1667.000 ;
        RECT 4.400 1641.160 2796.000 1642.560 ;
        RECT 4.000 1616.720 2796.000 1641.160 ;
        RECT 4.400 1615.320 2796.000 1616.720 ;
        RECT 4.000 1614.000 2796.000 1615.320 ;
        RECT 4.000 1612.600 2795.600 1614.000 ;
        RECT 4.000 1590.880 2796.000 1612.600 ;
        RECT 4.400 1589.480 2796.000 1590.880 ;
        RECT 4.000 1565.040 2796.000 1589.480 ;
        RECT 4.400 1563.640 2796.000 1565.040 ;
        RECT 4.000 1559.600 2796.000 1563.640 ;
        RECT 4.000 1558.200 2795.600 1559.600 ;
        RECT 4.000 1539.200 2796.000 1558.200 ;
        RECT 4.400 1537.800 2796.000 1539.200 ;
        RECT 4.000 1513.360 2796.000 1537.800 ;
        RECT 4.400 1511.960 2796.000 1513.360 ;
        RECT 4.000 1505.200 2796.000 1511.960 ;
        RECT 4.000 1503.800 2795.600 1505.200 ;
        RECT 4.000 1487.520 2796.000 1503.800 ;
        RECT 4.400 1486.120 2796.000 1487.520 ;
        RECT 4.000 1461.680 2796.000 1486.120 ;
        RECT 4.400 1460.280 2796.000 1461.680 ;
        RECT 4.000 1450.800 2796.000 1460.280 ;
        RECT 4.000 1449.400 2795.600 1450.800 ;
        RECT 4.000 1435.840 2796.000 1449.400 ;
        RECT 4.400 1434.440 2796.000 1435.840 ;
        RECT 4.000 1410.000 2796.000 1434.440 ;
        RECT 4.400 1408.600 2796.000 1410.000 ;
        RECT 4.000 1396.400 2796.000 1408.600 ;
        RECT 4.000 1395.000 2795.600 1396.400 ;
        RECT 4.000 1384.160 2796.000 1395.000 ;
        RECT 4.400 1382.760 2796.000 1384.160 ;
        RECT 4.000 1358.320 2796.000 1382.760 ;
        RECT 4.400 1356.920 2796.000 1358.320 ;
        RECT 4.000 1342.000 2796.000 1356.920 ;
        RECT 4.000 1340.600 2795.600 1342.000 ;
        RECT 4.000 1332.480 2796.000 1340.600 ;
        RECT 4.400 1331.080 2796.000 1332.480 ;
        RECT 4.000 1306.640 2796.000 1331.080 ;
        RECT 4.400 1305.240 2796.000 1306.640 ;
        RECT 4.000 1287.600 2796.000 1305.240 ;
        RECT 4.000 1286.200 2795.600 1287.600 ;
        RECT 4.000 1280.800 2796.000 1286.200 ;
        RECT 4.400 1279.400 2796.000 1280.800 ;
        RECT 4.000 1254.960 2796.000 1279.400 ;
        RECT 4.400 1253.560 2796.000 1254.960 ;
        RECT 4.000 1233.200 2796.000 1253.560 ;
        RECT 4.000 1231.800 2795.600 1233.200 ;
        RECT 4.000 1229.120 2796.000 1231.800 ;
        RECT 4.400 1227.720 2796.000 1229.120 ;
        RECT 4.000 1203.280 2796.000 1227.720 ;
        RECT 4.400 1201.880 2796.000 1203.280 ;
        RECT 4.000 1178.800 2796.000 1201.880 ;
        RECT 4.000 1177.440 2795.600 1178.800 ;
        RECT 4.400 1177.400 2795.600 1177.440 ;
        RECT 4.400 1176.040 2796.000 1177.400 ;
        RECT 4.000 1151.600 2796.000 1176.040 ;
        RECT 4.400 1150.200 2796.000 1151.600 ;
        RECT 4.000 1125.760 2796.000 1150.200 ;
        RECT 4.400 1124.400 2796.000 1125.760 ;
        RECT 4.400 1124.360 2795.600 1124.400 ;
        RECT 4.000 1123.000 2795.600 1124.360 ;
        RECT 4.000 1099.920 2796.000 1123.000 ;
        RECT 4.400 1098.520 2796.000 1099.920 ;
        RECT 4.000 1074.080 2796.000 1098.520 ;
        RECT 4.400 1072.680 2796.000 1074.080 ;
        RECT 4.000 1070.000 2796.000 1072.680 ;
        RECT 4.000 1068.600 2795.600 1070.000 ;
        RECT 4.000 1048.240 2796.000 1068.600 ;
        RECT 4.400 1046.840 2796.000 1048.240 ;
        RECT 4.000 1022.400 2796.000 1046.840 ;
        RECT 4.400 1021.000 2796.000 1022.400 ;
        RECT 4.000 1015.600 2796.000 1021.000 ;
        RECT 4.000 1014.200 2795.600 1015.600 ;
        RECT 4.000 996.560 2796.000 1014.200 ;
        RECT 4.400 995.160 2796.000 996.560 ;
        RECT 4.000 970.720 2796.000 995.160 ;
        RECT 4.400 969.320 2796.000 970.720 ;
        RECT 4.000 961.200 2796.000 969.320 ;
        RECT 4.000 959.800 2795.600 961.200 ;
        RECT 4.000 944.880 2796.000 959.800 ;
        RECT 4.400 943.480 2796.000 944.880 ;
        RECT 4.000 919.040 2796.000 943.480 ;
        RECT 4.400 917.640 2796.000 919.040 ;
        RECT 4.000 906.800 2796.000 917.640 ;
        RECT 4.000 905.400 2795.600 906.800 ;
        RECT 4.000 893.200 2796.000 905.400 ;
        RECT 4.400 891.800 2796.000 893.200 ;
        RECT 4.000 867.360 2796.000 891.800 ;
        RECT 4.400 865.960 2796.000 867.360 ;
        RECT 4.000 852.400 2796.000 865.960 ;
        RECT 4.000 851.000 2795.600 852.400 ;
        RECT 4.000 841.520 2796.000 851.000 ;
        RECT 4.400 840.120 2796.000 841.520 ;
        RECT 4.000 815.680 2796.000 840.120 ;
        RECT 4.400 814.280 2796.000 815.680 ;
        RECT 4.000 798.000 2796.000 814.280 ;
        RECT 4.000 796.600 2795.600 798.000 ;
        RECT 4.000 789.840 2796.000 796.600 ;
        RECT 4.400 788.440 2796.000 789.840 ;
        RECT 4.000 764.000 2796.000 788.440 ;
        RECT 4.400 762.600 2796.000 764.000 ;
        RECT 4.000 743.600 2796.000 762.600 ;
        RECT 4.000 742.200 2795.600 743.600 ;
        RECT 4.000 738.160 2796.000 742.200 ;
        RECT 4.400 736.760 2796.000 738.160 ;
        RECT 4.000 712.320 2796.000 736.760 ;
        RECT 4.400 710.920 2796.000 712.320 ;
        RECT 4.000 689.200 2796.000 710.920 ;
        RECT 4.000 687.800 2795.600 689.200 ;
        RECT 4.000 686.480 2796.000 687.800 ;
        RECT 4.400 685.080 2796.000 686.480 ;
        RECT 4.000 660.640 2796.000 685.080 ;
        RECT 4.400 659.240 2796.000 660.640 ;
        RECT 4.000 634.800 2796.000 659.240 ;
        RECT 4.400 633.400 2795.600 634.800 ;
        RECT 4.000 608.960 2796.000 633.400 ;
        RECT 4.400 607.560 2796.000 608.960 ;
        RECT 4.000 583.120 2796.000 607.560 ;
        RECT 4.400 581.720 2796.000 583.120 ;
        RECT 4.000 580.400 2796.000 581.720 ;
        RECT 4.000 579.000 2795.600 580.400 ;
        RECT 4.000 557.280 2796.000 579.000 ;
        RECT 4.400 555.880 2796.000 557.280 ;
        RECT 4.000 531.440 2796.000 555.880 ;
        RECT 4.400 530.040 2796.000 531.440 ;
        RECT 4.000 526.000 2796.000 530.040 ;
        RECT 4.000 524.600 2795.600 526.000 ;
        RECT 4.000 505.600 2796.000 524.600 ;
        RECT 4.400 504.200 2796.000 505.600 ;
        RECT 4.000 479.760 2796.000 504.200 ;
        RECT 4.400 478.360 2796.000 479.760 ;
        RECT 4.000 471.600 2796.000 478.360 ;
        RECT 4.000 470.200 2795.600 471.600 ;
        RECT 4.000 453.920 2796.000 470.200 ;
        RECT 4.400 452.520 2796.000 453.920 ;
        RECT 4.000 428.080 2796.000 452.520 ;
        RECT 4.400 426.680 2796.000 428.080 ;
        RECT 4.000 417.200 2796.000 426.680 ;
        RECT 4.000 415.800 2795.600 417.200 ;
        RECT 4.000 402.240 2796.000 415.800 ;
        RECT 4.400 400.840 2796.000 402.240 ;
        RECT 4.000 376.400 2796.000 400.840 ;
        RECT 4.400 375.000 2796.000 376.400 ;
        RECT 4.000 362.800 2796.000 375.000 ;
        RECT 4.000 361.400 2795.600 362.800 ;
        RECT 4.000 350.560 2796.000 361.400 ;
        RECT 4.400 349.160 2796.000 350.560 ;
        RECT 4.000 324.720 2796.000 349.160 ;
        RECT 4.400 323.320 2796.000 324.720 ;
        RECT 4.000 308.400 2796.000 323.320 ;
        RECT 4.000 307.000 2795.600 308.400 ;
        RECT 4.000 298.880 2796.000 307.000 ;
        RECT 4.400 297.480 2796.000 298.880 ;
        RECT 4.000 273.040 2796.000 297.480 ;
        RECT 4.400 271.640 2796.000 273.040 ;
        RECT 4.000 254.000 2796.000 271.640 ;
        RECT 4.000 252.600 2795.600 254.000 ;
        RECT 4.000 247.200 2796.000 252.600 ;
        RECT 4.400 245.800 2796.000 247.200 ;
        RECT 4.000 221.360 2796.000 245.800 ;
        RECT 4.400 219.960 2796.000 221.360 ;
        RECT 4.000 199.600 2796.000 219.960 ;
        RECT 4.000 198.200 2795.600 199.600 ;
        RECT 4.000 195.520 2796.000 198.200 ;
        RECT 4.400 194.120 2796.000 195.520 ;
        RECT 4.000 169.680 2796.000 194.120 ;
        RECT 4.400 168.280 2796.000 169.680 ;
        RECT 4.000 145.200 2796.000 168.280 ;
        RECT 4.000 143.840 2795.600 145.200 ;
        RECT 4.400 143.800 2795.600 143.840 ;
        RECT 4.400 142.440 2796.000 143.800 ;
        RECT 4.000 118.000 2796.000 142.440 ;
        RECT 4.400 116.600 2796.000 118.000 ;
        RECT 4.000 92.160 2796.000 116.600 ;
        RECT 4.400 90.800 2796.000 92.160 ;
        RECT 4.400 90.760 2795.600 90.800 ;
        RECT 4.000 89.400 2795.600 90.760 ;
        RECT 4.000 66.320 2796.000 89.400 ;
        RECT 4.400 64.920 2796.000 66.320 ;
        RECT 4.000 40.480 2796.000 64.920 ;
        RECT 4.400 39.080 2796.000 40.480 ;
        RECT 4.000 36.400 2796.000 39.080 ;
        RECT 4.000 35.000 2795.600 36.400 ;
        RECT 4.000 14.640 2796.000 35.000 ;
        RECT 4.400 13.240 2796.000 14.640 ;
        RECT 4.000 2.895 2796.000 13.240 ;
      LAYER met4 ;
        RECT 868.775 10.240 942.240 1557.025 ;
        RECT 944.640 10.240 1019.040 1557.025 ;
        RECT 1021.440 10.240 1095.840 1557.025 ;
        RECT 1098.240 10.240 1172.640 1557.025 ;
        RECT 1175.040 10.240 1249.440 1557.025 ;
        RECT 1251.840 10.240 1326.240 1557.025 ;
        RECT 1328.640 10.240 1403.040 1557.025 ;
        RECT 1405.440 10.240 1479.840 1557.025 ;
        RECT 1482.240 10.240 1556.640 1557.025 ;
        RECT 1559.040 10.240 1632.705 1557.025 ;
        RECT 868.775 3.575 1632.705 10.240 ;
  END
END picorv32
END LIBRARY

